module ceshi #(
    parameters
) (
    input clk ,
    input rst ,
    output  led 
);


    
endmodule